// fixedDSP.v

// Generated using ACDS version 19.1 240

`timescale 1 ps / 1 ps
module fixedDSP (
		input  wire [17:0] ay,      //      ay.ay
		input  wire [17:0] by,      //      by.by
		input  wire [17:0] ax,      //      ax.ax
		input  wire [17:0] bx,      //      bx.bx
		output wire [36:0] resulta, // resulta.resulta
		output wire [36:0] resultb  // resultb.resultb
	);

	fixedDSP_altera_c10gx_native_fixed_point_dsp_191_g2gyhoq c10gx_native_fixed_point_dsp_0 (
		.ay      (ay),      //   input,  width = 18,      ay.ay
		.by      (by),      //   input,  width = 18,      by.by
		.ax      (ax),      //   input,  width = 18,      ax.ax
		.bx      (bx),      //   input,  width = 18,      bx.bx
		.resulta (resulta), //  output,  width = 37, resulta.resulta
		.resultb (resultb)  //  output,  width = 37, resultb.resultb
	);

endmodule
