module issp (
		output wire [17:0] source, // sources.source
		input  wire [99:0] probe   //  probes.probe
	);
endmodule

