module fixedDSP (
		input  wire [17:0] ay,      //      ay.ay
		input  wire [17:0] by,      //      by.by
		input  wire [17:0] ax,      //      ax.ax
		input  wire [17:0] bx,      //      bx.bx
		output wire [63:0] resulta  // resulta.resulta
	);
endmodule

