module parallel_add (
		input  wire [15:0] data0x, //  parallel_add_input.data0x
		input  wire [15:0] data1x, //                    .data1x
		input  wire [15:0] data2x, //                    .data2x
		input  wire [15:0] data3x, //                    .data3x
		input  wire [15:0] data4x, //                    .data4x
		output wire [18:0] result  // parallel_add_output.result
	);
endmodule

