// paral_add.v

// Generated using ACDS version 19.1 240

`timescale 1 ps / 1 ps
module paral_add (
		input  wire [15:0] data0x, //  parallel_add_input.data0x
		input  wire [15:0] data1x, //                    .data1x
		input  wire [15:0] data2x, //                    .data2x
		input  wire [15:0] data3x, //                    .data3x
		input  wire [15:0] data4x, //                    .data4x
		output wire [18:0] result  // parallel_add_output.result
	);

	paral_add_parallel_add_191_u2agy2i parallel_add_0 (
		.data0x (data0x), //   input,  width = 16,  parallel_add_input.data0x
		.data1x (data1x), //   input,  width = 16,                    .data1x
		.data2x (data2x), //   input,  width = 16,                    .data2x
		.data3x (data3x), //   input,  width = 16,                    .data3x
		.data4x (data4x), //   input,  width = 16,                    .data4x
		.result (result)  //  output,  width = 19, parallel_add_output.result
	);

endmodule
