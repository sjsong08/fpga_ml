module issp2 (
		output wire [0:0]   source, // sources.source
		input  wire [437:0] probe   //  probes.probe
	);
endmodule

