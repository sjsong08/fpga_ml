// bram_24.v

// Generated using ACDS version 18.1 222

`timescale 1 ps / 1 ps
module bram_24 (
		input  wire [23:0] data,    //    data.datain
		output wire [23:0] q,       //       q.dataout
		input  wire [10:0] address, // address.address
		input  wire        wren,    //    wren.wren
		input  wire        clock,   //   clock.clk
		input  wire        rden     //    rden.rden
	);

	bram_24_ram_1port_181_w7eesfi ram_1port_0 (
		.data    (data),    //   input,  width = 24,    data.datain
		.q       (q),       //  output,  width = 24,       q.dataout
		.address (address), //   input,  width = 11, address.address
		.wren    (wren),    //   input,   width = 1,    wren.wren
		.clock   (clock),   //   input,   width = 1,   clock.clk
		.rden    (rden)     //   input,   width = 1,    rden.rden
	);

endmodule
