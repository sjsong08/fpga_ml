module issp (
		output wire [3:0]  source, // sources.source
		input  wire [47:0] probe   //  probes.probe
	);
endmodule

