module issp (
		output wire [2:0]   source, // sources.source
		input  wire [351:0] probe   //  probes.probe
	);
endmodule

