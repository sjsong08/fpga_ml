module para_add (
		input  wire [18:0] data0x, //  parallel_add_input.data0x
		input  wire [18:0] data1x, //                    .data1x
		input  wire [18:0] data2x, //                    .data2x
		output wire [20:0] result  // parallel_add_output.result
	);
endmodule

