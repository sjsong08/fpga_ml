module stp (
		input  wire [79:0] acq_data_in,    //     tap.acq_data_in
		input  wire [2:0]  acq_trigger_in, //        .acq_trigger_in
		input  wire        acq_clk         // acq_clk.clk
	);
endmodule

