module stp (
		input  wire [9:0] acq_data_in,    //     tap.acq_data_in
		input  wire [0:0] acq_trigger_in, //        .acq_trigger_in
		input  wire       acq_clk         // acq_clk.clk
	);
endmodule

